            logic [7:0] uart_status;            logic [7:0] uart_send_byte;            logic [7:0] uart_rcvd_byte;            logic [7:0] uart_cfg;