module if(
    input               clk,
    input        [31:0] i_data_in,
    input        [31:0] i_addr,
    output logic [31:0] i_addr,
    output logic [31:0] i_data_out
);
    logic [31:0] prev_data;
    always @(posedge clk) begin
    end

endmodule
