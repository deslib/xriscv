module tb_soc;
endmodule
